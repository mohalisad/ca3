`timescale 1ns/1ns
module instructreg(input[12:0] in,input rst,output reg[7:0] out);
	reg[7:0]r[0:8191];
	always@(in,rst)begin
		r[0]<=8'b01000011;
		r[1]<=8'b11101000;
		r[2]<=8'b10010110;
		r[3]<=8'b01000011;
		r[4]<=8'b11101001;
		r[5]<=8'b10010110;
		r[6]<=8'b01000011;
		r[7]<=8'b11101010;
		r[8]<=8'b10010110;
		r[9]<=8'b01000011;
		r[10]<=8'b11101011;
		r[11]<=8'b10010110;
		r[12]<=8'b01000011;
		r[13]<=8'b11101100;
		r[14]<=8'b10010110;
		r[15]<=8'b01000011;
		r[16]<=8'b11101101;
		r[17]<=8'b10010110;
		r[18]<=8'b01000011;
		r[19]<=8'b11101110;
		r[20]<=8'b10010110;
		r[21]<=8'b01000011;
		r[22]<=8'b11101111;
		r[23]<=8'b10010110;
		r[24]<=8'b01000011;
		r[25]<=8'b11110000;
		r[26]<=8'b10010110;
		r[27]<=8'b01000011;
		r[28]<=8'b11110001;
		r[29]<=8'b10010110;

		r[30]<=8'b00100111;
		r[31]<=8'b11010000;

		r[32]<=8'b11101000;

		r[33]<=8'b00100111;
		r[34]<=8'b11010001;
		r[8191]<=8'b11100000;
		if(rst)
			out<=0;
		else
			out<=r[in];
	end
endmodule
